module Garnet_TB (
                  input         clk,
                  input         reset,
                  output        GC_interrupt,
                  input [12:0]  GC_ARADDR,
                  output        GC_ARREADY,
                  input         GC_ARVALID,
                  input [12:0]  GC_AWADDR,
                  output        GC_AWREADY,
                  input         GC_AWVALID,
                  output [31:0] GC_RDATA,
                  input         GC_RREADY,
                  output [1:0]  GC_RRESP,
                  output        GC_RVALID,
                  input [31:0]  GC_WDATA,
                  output        GC_WREADY,
                  input         GC_WVALID,
                  input [3:0]   GC_WSTRB,
                  output        GC_BVALID,
                  input         GC_BREADY,
                  output [1:0]  GC_BRESP,
                  input         JTAG_TCK,
                  input         JTAG_TDI,
                  output        JTAG_TDO,
                  input         JTAG_TMS,
                  input         JTAG_TRSTn,
                  input [31:0]  GB_rd_addr,
                  output [63:0] GB_rd_data,
                  output        GB_rd_data_valid,
                  input         GB_rd_en,
                  input [31:0]  GB_wr_addr,
                  input [63:0]  GB_wr_data,
                  input         GB_wr_en,
                  input [7:0]   GB_wr_strb,
                  input         TB_monitor_power
                  );

   Garnet DUT (.clk_in(clk),
               .reset_in(reset),
               .axi4_slave_araddr(GC_ARADDR),
               .axi4_slave_arready(GC_ARREADY),
               .axi4_slave_arvalid(GC_ARVALID),
               .axi4_slave_awaddr(GC_AWADDR),
               .axi4_slave_awready(GC_AWREADY),
               .axi4_slave_awvalid(GC_AWVALID),
               .axi4_slave_bready(GC_BREADY),
               .axi4_slave_bresp(GC_BRESP),
               .axi4_slave_bvalid(GC_BVALID),
               .axi4_slave_rdata(GC_RDATA),
               .axi4_slave_rready(GC_RREADY),
               .axi4_slave_rresp(GC_RRESP),
               .axi4_slave_rvalid(GC_RVALID),
               .axi4_slave_wdata(GC_WDATA),
               .axi4_slave_wready(GC_WREADY),
               .axi4_slave_wvalid(GC_WVALID),
               .interrupt(GC_interrupt),
               .jtag_tck(JTAG_TCK),
               .jtag_tdi(JTAG_TDI),
               .jtag_tdo(JTAG_TDO),
               .jtag_tms(JTAG_TMS),
               .jtag_trst_n(JTAG_TRSTn),
               .proc_packet_rd_addr(GB_rd_addr),
               .proc_packet_rd_data(GB_rd_data),
               .proc_packet_rd_data_valid(GB_rd_data_valid),
               .proc_packet_rd_en(GB_rd_en),
               .proc_packet_wr_addr(GB_wr_addr),
               .proc_packet_wr_data(GB_wr_data),
               .proc_packet_wr_en(GB_wr_en),
               .proc_packet_wr_strb(GB_wr_strb)
               );

endmodule // Garnet_TB
