module Garnet_TB (
                  input         clk,
                  input         reset,
                  output        GC_interrupt,
                  input [11:0]  GC_ARADDR,
                  output        GC_ARREADY,
                  input         GC_ARVALID,
                  input [11:0]  GC_AWADDR,
                  output        GC_AWREADY,
                  input         GC_AWVALID,
                  output [31:0] GC_RDATA,
                  input         GC_RREADY,
                  output [1:0]  GC_RRESP,
                  output        GC_RVALID,
                  input [31:0]  GC_WDATA,
                  output        GC_WREADY,
                  input         GC_WVALID,
                  input [3:0]   GC_WSTRB,
                  output        GC_BVALID,
                  input         GC_BREADY,
                  output        GC_BRESP,
                  input         JTAG_TCK,
                  input         JTAG_TDI,
                  output        JTAG_TDO,
                  input         JTAG_TMS,
                  input         JTAG_TRSTn,
                  input [31:0]  GB_rd_addr,
                  output [63:0] GB_rd_data,
                  input         GB_rd_en,
                  input [31:0]  GB_wr_addr,
                  input [63:0]  GB_wr_data,
                  input [7:0]   GB_wr_strb,
                  input         TB_monitor_power
                  );

   assign GC_BVALID = 1;
   assign GC_BRESP = 0;

   Garnet DUT (.clk_in(clk),
               .reset_in(reset),
               .axi4_ctrl_araddr(GC_ARADDR),
               .axi4_ctrl_arready(GC_ARREADY),
               .axi4_ctrl_arvalid(GC_ARVALID),
               .axi4_ctrl_awaddr(GC_AWADDR),
               .axi4_ctrl_awready(GC_AWREADY),
               .axi4_ctrl_awvalid(GC_AWVALID),
               .axi4_ctrl_rdata(GC_RDATA),
               .axi4_ctrl_rready(GC_RREADY),
               .axi4_ctrl_rresp(GC_RRESP),
               .axi4_ctrl_rvalid(GC_RVALID),
               .axi4_ctrl_wdata(GC_WDATA),
               .axi4_ctrl_wready(GC_WREADY),
               .axi4_ctrl_wvalid(GC_WVALID),
               .axi4_ctrl_interrupt(GC_interrupt),
               .jtag_tck(JTAG_TCK),
               .jtag_tdi(JTAG_TDI),
               .jtag_tdo(JTAG_TDO),
               .jtag_tms(JTAG_TMS),
               .jtag_trst_n(JTAG_TRSTn),
               .soc_data_rd_addr(GB_rd_addr),
               .soc_data_rd_data(GB_rd_data),
               .soc_data_rd_en(GB_rd_en),
               .soc_data_wr_addr(GB_wr_addr),
               .soc_data_wr_data(GB_wr_data),
               .soc_data_wr_strb(GB_wr_strb)
               );

endmodule // Garnet_TB
